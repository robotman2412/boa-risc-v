
// Copyright © 2024, Julian Scheffers, see LICENSE for more information

`timescale 1ns/1ps



module mmio_vga_periph(
    // VGA core clock.
    input  logic    vga_clk,
    // Memory bus clock.
    input  logic    mem_clk,
);
endmodule
